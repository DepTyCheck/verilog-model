// Seed: 18199170163325466416,2426731264514140405

module zh
  (output logic [2:2] nebhihq, output uwire bqj, output logic ayneqzd, output logic [4:3] blfhjlbbph, input bit [1:0] hyq);
  
  
  and xuqytvefhf(pqxmjgo, nebhihq, ayneqzd);
  
  not yuiohpctmh(ayneqzd, hkr);
  
  not aamvrptl(nebhihq, hqcrpoga);
  
  
  // Top inputs -> top outputs assigns
  
  // Assigns
  assign hqcrpoga = 'b1;
  assign hqcrpoga = 'bx;
  assign bqj = 'b1;
  assign blfhjlbbph = 'b1z;
  assign pqxmjgo = 'bz;
  assign pqxmjgo = 'bz;
endmodule: zh



// Seed after: 11453228651617964993,2426731264514140405
