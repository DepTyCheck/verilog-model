// Seed: 11453228651617964993,2426731264514140405

module fzasj
  (output real plufmmppl [0:3][0:4], output int gfezbggpe, output bit [2:3][4:2] gwxcoakrzk, output bit [2:1] spuvn);
  
  
  not zk(gwxcoakrzk, gwxcoakrzk);
  // warning: implicit conversion of port connection expands from 1 to 6 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic gwxcoakrzk -> bit [2:3][4:2] gwxcoakrzk
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:3][4:2] gwxcoakrzk -> logic gwxcoakrzk
  
  not yfhwyau(jholzoq, gp);
  
  nand ake(sfi, zyjksdtagv, jholzoq);
  
  or m(spuvn, hjpy, spuvn);
  // warning: implicit conversion of port connection expands from 1 to 2 bits
  // warning: implicit conversion changes possible bit states from 4-state to 2-state
  //   logic spuvn -> bit [2:1] spuvn
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:1] spuvn -> logic spuvn
  
  
  // Top inputs -> top outputs assigns
  
  // Assigns
  assign hjpy = 'bz;
  assign zyjksdtagv = 'b0;
  assign gp = 'b0;
  assign gfezbggpe = 'b0;
  assign plufmmppl = '{'{'b1,'b0,'b1,'bx,'bx},'{'bz,'bz,'b1,'b1,'b0},'{'b1,'bx,'bx,'bx,'b1},'{'b0,'bz,'bz,'bx,'b0}};
  assign jholzoq = 'b1;
  assign sfi = 'bz;
endmodule: fzasj

module etvas
  ();
  
  
  not qcglhthwsu(uniktucuj, xkveoe);
  
  and yupqw(d, jgazddhls, ofbgbhkoo);
  
  not gdybviu(ofbgbhkoo, xcyfoyomq);
  
  
  // Top inputs -> top outputs assigns
  
  // Assigns
  assign d = 'bz;
endmodule: etvas

module v
  (output logic [2:3] f [3:1], output logic [1:2] o [4:0]);
  
  real xnyvbyx [0:3][0:4];
  
  fzasj erus(.plufmmppl(xnyvbyx), .gfezbggpe(nyla), .gwxcoakrzk(zbyunv), .spuvn(zqwt));
  // warning: implicit conversion of port connection truncates from 32 to 1 bits
  // warning: implicit conversion changes signedness from signed to unsigned
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   int gfezbggpe -> wire nyla
  //
  // warning: implicit conversion of port connection truncates from 6 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:3][4:2] gwxcoakrzk -> wire zbyunv
  //
  // warning: implicit conversion of port connection truncates from 2 to 1 bits
  // warning: implicit conversion changes possible bit states from 2-state to 4-state
  //   bit [2:1] spuvn -> wire zqwt
  
  etvas ncn();
  
  not jxtvshncq(lkxtjzty, nyla);
  
  
  // Top inputs -> top outputs assigns
  
  // Assigns
  assign nyla = 'bx;
endmodule: v



// Seed after: 5123120746938755423,2426731264514140405
