entity helloworld is
end helloworld;

architecture behaviour of helloworld is
begin
end behaviour;

entity lmao is
end lmao;

architecture behaviour2 of lmao is
begin
end behaviour2;
