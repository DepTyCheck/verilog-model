// Seed: 18347911916735053405,2426731264514140405

module zbjft
  (output real hftsz [2:1], output bit rhqocjml [1:1], output int dyhck);
  
  
  xor bauagpzq(mmchqmwvv, ctophjw, vh);
  
  
  // Top inputs -> top outputs assigns
  
  // Assigns
  assign vh = 'bx;
  assign ctophjw = 'b0;
  assign hftsz = '{'bx,'bx};
  assign mmchqmwvv = 'b0;
  assign mmchqmwvv = 'b1;
endmodule: zbjft

module agxj
  ( output integer uvujoem [1:0]
  , output wire cgpe [4:1]
  , output logic pwhnwwmffv [4:3]
  , output bit [2:1][3:3] w
  , input real cesmyxprke
  , input logic [2:3] ajkuhiz
  , input bit [4:0] yjjdnwp
  , input uwire ue
  );
  
  
  
  // Top inputs -> top outputs assigns
  
  // Assigns
  assign w = 'b10;
  assign pwhnwwmffv = '{'b0,'bx};
  assign uvujoem = '{'b0,'b0};
  assign cgpe = '{'b0,'b0,'b0,'b0};
endmodule: agxj



// Seed after: 12155394080032148100,2426731264514140405
